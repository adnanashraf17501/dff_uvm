module DUT(intif.dut inf);
df vcode(.clk(inf.clk),.rst(inf.rst),.d(inf.d),.q(inf.q));
endmodule
